`define ST_IDLE 3'd0
`define ST_LOAD_A 3'd1
`define ST_LOAD_B 3'd2
`define ST_LOAD_OP 3'd3
`define ST_DONE_A  3'd5
`define ST_DONE_B  3'd6
`define ST_DONE_OP 3'd7