`define OP_ADD 4'd0
`define OP_SUB 4'd1
`define OP_AND 4'd2
`define OP_OR  4'd3
`define OP_XOR 4'd4
`define OP_PASS_A 4'd5
`define OP_PASS_B 4'd6
`define OP_SHL_A  4'd7
`define OP_SHR_A  4'd8
`define OP_MOVE_REG_XA 4'd9 // move a to x
`define OP_MOVE_REG_AX 4'd10 // move x to a
`define OP_INC_REG_A 4'd11
`define OP_DEC_REG_A 4'd12