`define OP_ADD 5'd0
`define OP_SUB 5'd1
`define OP_AND 5'd2
`define OP_OR 5'd3
`define OP_XOR 5'd4
`define OP_PASS_A 5'd5
`define OP_PASS_B 5'd6
`define OP_SHL_A 5'd7
`define OP_SHR_A 5'd8
`define OP_MOVE_REG_XA 5'd9 // move a to x
`define OP_MOVE_REG_AX 5'd10 // move x to a
`define OP_INC_REG_A 5'd11
`define OP_DEC_REG_A 5'd12
`define OP_NOT_A 5'd13
`define OP_NEG_A 5'd14
`define OP_CLR_A 5'd15
`define OP_MAX 5'd16
`define OP_MIN 5'd17
`define OP_ABS_A 5'd18